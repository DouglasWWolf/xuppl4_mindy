
//================================================================================================
//    Date         Version  Who  Changes
// -----------------------------------------------------------------------------------------------
// 22-Feb-2024       1.0.0  DWW  Initial creation
//================================================================================================
localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 0;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0;

localparam VERSION_MONTH = 2;
localparam VERSION_DAY   = 22;
localparam VERSION_YEAR  = 2024;
