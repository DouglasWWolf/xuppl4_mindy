
//================================================================================================
//    Date         Version  Who  Changes
// -----------------------------------------------------------------------------------------------
// 22-Feb-2024       1.0.0  DWW  Initial creation
//
// 24-Mar-2024       2.0.0  DWW  Added the abm-manager
//================================================================================================
localparam VERSION_MAJOR = 2;
localparam VERSION_MINOR = 0;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0;

localparam VERSION_MONTH = 3;
localparam VERSION_DAY   = 24;
localparam VERSION_YEAR  = 2024;
